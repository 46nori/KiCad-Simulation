.MODEL M_1N4148 D (
+IS       = 5.29582e-09    
+RS       = 0.373588       N        = 1.68058        
+BV       = 110            IBV      = 5e-05          CJO      = 1.15e-12       
+VJ       = 0.737407       MJ       = 0.020644       FC       = 0.5            
+AF       = 1              XTI      = 3.80469        
+EG       = 1.10578        TRS1     = 1.69802e-06    TRS2     = 0              
+KF       = 0              TNOM     = 27             TT       = 5.19183e-10 )